//2.-CONTROL DE MOTOR A PASOS:
//Modulo que usa el divisor de reloj para prender y apagar las 2 bobinas A y B del motor a pasos bipolar
//de tipo NEMA 17, este motor cuenta con un controlador A4988 y a traves de sus pines STEP Y DIR se puede 
//controlar su movimiento y sentido de giro, cada vez que el pin STEP reciba un pulso, dara un paso, la 
//mayoria de motores bipolares dan pasos 200 pasos para dar una vuelta completa, osea que dan un giro de 
//1.8 grados, algunos dan giros de 400 pasos, osea 0.9 grados de rotacion por paso. 
//En el motor bipolar se cuenta con 5 secuencias de pasos principales: Paso completo, medio paso, 1/4 de 
//paso, 1/8 de paso y 1/16 de paso, mientras mas se disminuya el paso, mejor sera la precision de su 
//movimiento, pero su torque se reducira proporcionalmente, el torque maximo del motor se alcanza en el 
//paso completo, donde aguanta hasta 4kg de peso en una carga.

module controlPasosMotor(
	 input direccionGiro,
	 input [2:0] selectPaso,
	 //Se pueden elegir 5 opciones de pasos: Paso Completo, 1/2 paso, 1/4 de paso, 1/8 de paso y 1/16 de paso.
	 //Mientras sea menor el paso, mayor sera su precision, pero se reduce su torque de forma proporcional.
    output reg [2:0] MS, //Las salidas usadas dentro de un condicional o bucle se declaran como reg.
	 output reg [2:0] ledMS,
	 output reg DIR,
	 output reg ledDireccion
    );
	
	//always@() sirve para hacer operaciones matematicas, condicionales o bucles, dentro de su parentesis se 
	//deben poner las entradas que usara y ademas tiene su propio begin y end.
	always@(direccionGiro, selectPaso)
	begin
		//CONDICIONAL CASE: Se usa para evaluar los diferentes valores de la variable que tenga en su 
		//parentesis y asignar una salida correspondiente a cada caso.
		case(selectPaso)
			//Con los 3 pines MS1, MS2 y MS3 de Micro Stepping (MS), se establece el tipo de paso del motor para
			//lograr una mayor precision o torque, se elige una de las siguientes opciones:
			//							MS1	MS2	MS3	
			//Paso Completo = 	 0		 0		 0
			//Paso Medio = 	    1		 0		 0
			//1/4 de Paso = 	    0		 1		 0
			//1/8 de Paso = 	    1		 1		 0
			//1/16 de Paso = 	    1		 1		 1
			//Mientras mas se reduzca el paso, mayor es la resolucion de la precision en su movimiento, pero el 
			//torque se reduce proporcionalmente:
			//# Pasos 1 vuelta paso completo = 200 [pasos/revolucion]
			//# Pasos 1 vuelta cualquier otro paso = # Pasos 1 vuelta paso completo * 1/division de paso
			//# Pasos 1 vuelta de 1/4 de paso = 200 * 1/(1/4) = 200 * 4 = 800 [pasos/revolucion]
			3'b000 : begin MS = 3'b000; ledMS = 3'b000; end		//Paso completo.
			3'b001 : begin MS = 3'b100; ledMS = 3'b100; end		//1/2 Paso.
			3'b010 : begin MS = 3'b010; ledMS = 3'b010; end		//1/4 de Paso.
			3'b011 : begin MS = 3'b110; ledMS = 3'b110; end		//1/8 de Paso.
			3'b100 : begin MS = 3'b111; ledMS = 3'b111; end		//1/16 de Paso.
			//Si quiero que se ejecute algo cuando no se cumpla ninguna de las dos condiciones anteriores uso 
			//default.
			default : begin MS = 3'b000; ledMS = 3'b000; end 	//Motor a pasos bipolar con paso completo.
		endcase
		if(direccionGiro == 1'b1) begin 
			DIR = 1'b1;	//DIR = 1; Giro del motor en sentido de las manecillas del reloj (derecha).
			ledDireccion = 1'b1;
		end else begin
			DIR = 1'b0;	//DIR = 0; Giro del motor en sentido contrario de las manecillas del reloj (izquierda).
			ledDireccion = 1'b0;
		end
	end
endmodule
